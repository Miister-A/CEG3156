-- nBit_cla4_adder

-- n must be a multiple of 4

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

entity nBit_cla4_adder is
	generic ( n : positive := 4 );
	port(
		a, b : in std_logic_vector(n-1 downto 0);
		c_in : in std_logic;
		sum : out std_logic_vector(n-1 downto 0);
		c_out, overflow : out std_logic);
end nBit_cla4_adder;

architecture structural of nBit_cla4_adder is

component cla4_adder is
	port(
		a, b : in std_logic_vector(3 downto 0);
		c_in : in std_logic;
		sum : out std_logic_vector(3 downto 0);
		c_ovfl, c_out : out std_logic);
end component;
		
signal c_in_mid, c_out_mid, c_ovfl_mid : std_logic_vector(n/4 downto 0);

begin
	assert (n mod 4 = 0) report "n must be a multiple of 4 for use in nBit_cla4_adder" severity FAILURE;

	c_in_mid(0) <= c_in;
	c_in_mid(n/4 downto 1) <= c_out_mid((n/4)-1 downto 0);
	c_out <= c_out_mid((n/4)-1);

	loop0: for i in 0 to ((n/4)-1) generate
		cla4_adder_inst : cla4_adder
			port map (a((i*4 + 3) downto (i*4)), 
						 b((i*4 + 3) downto (i*4)), 
						 c_in_mid(i), 
						 sum((i*4 + 3) downto (i*4)), 
						 c_ovfl_mid(i), 			-- only the last overflow bit is used
						 c_out_mid(i));
						 
	end generate;
	
	
	overflow <= c_in_mid((n/4)-1) xor c_ovfl_mid((n/4)-1);

end structural;